`ifndef __EXEC_CORE_PKG_SV__
`define __EXEC_CORE_PKG_SV__

`timescale 1ns / 1ns

`include "uvm_macros.svh"

package exec_core_pkg;

	import uvm_pkg::*;

	// `include "exec_core_transaction.sv"
	// `include "exec_core_driver.sv"
	// `include "exec_core_monitor.sv"
	// `include "exec_core_agent.sv"
	// `include "exec_core_sequence.sv"
	// `include "exec_core_scoreboard.sv"
	// `include "register_file_probe_if.sv"
	// `include "register_file_probe_config.sv"
	// `include "register_file_probe.sv"
	// `include "exec_core_env.sv"
//	`include "exec_core_tests.sv"

endpackage: exec_core_pkg

`endif

`timescale 1ns / 1ns

class exec_core_sequence extends uvm_sequence #(exec_core_transaction);

	`uvm_object_utils(exec_core_sequence)

	function new (string name = "");
		super.new(name);
	endfunction

	task body;
		`uvm_info(get_type_name(), "Sequence start", UVM_MEDIUM)
		// Perform an initial RESET to clean up the cpu state
		`uvm_do_with(req, { req.cmd == CMD_RESET; })
		repeat(2)
		begin
			`uvm_do_with(req, { req.cmd == CMD_ADDI; })
			// `uvm_do(req)
		end
	endtask: body

endclass: exec_core_sequence
